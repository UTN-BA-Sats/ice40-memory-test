`include "memory.v"

module MemorySet(
    input clk,
    input reset,
    input [7:0] addr,
    input [19:0] cs,
    input read_byte_sel,
    input rw,
    input [15:0] i_data_word,
    output [7:0] o_data_byte
);

Memory memory_inst0(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[0]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst0.INIT_0 = 256'hedc176b13db130c855f9dd712ec6ddfe9976709a3d2a4d634de00f2d629fe86d;
defparam memory_inst0.INIT_1 = 256'h52dcb7b6b965f7058504f603525440be0f1952b0b46df6a32cabb007d95790bb;
defparam memory_inst0.INIT_2 = 256'h52fd4ec397e2f42c262eaaeb40773d8d89361865937ce8e39041286f7b07fbab;
defparam memory_inst0.INIT_3 = 256'hd8d7e5f4ab378a574e6b6a17cf8921c18e603c7b7836eb575d38e5f37f9b42ee;
defparam memory_inst0.INIT_4 = 256'h619caf9dca8add41b1d9cef1ed570d20c0a86ad30b6a84cd762da2722c92abf3;
defparam memory_inst0.INIT_5 = 256'h3368e70cca148a6e3a3f5445aacc7834e15c17f457cba183bfbbe3da73c25993;
defparam memory_inst0.INIT_6 = 256'h4f03d9c99225d03454eac518a9830a1e53326105e6ed942a72445e6a760c920e;
defparam memory_inst0.INIT_7 = 256'hdd8d647842f541b19e3415d1838b6794446b577863cd22e3e88dccdaf2446c7f;
defparam memory_inst0.INIT_8 = 256'he2902e0eb2647eeff7d4a6a6b057144a430de280d0c9f3e0038c46935470df68;
defparam memory_inst0.INIT_9 = 256'he6a3de90ec643ddea0e4798a9b6de728593bb1cd4d8c1f01b8499014b69bbea7;
defparam memory_inst0.INIT_A = 256'h01ea8716c1abb00f7b3ef228360ff85ba4b63a5eb955690955e2f217b7b6e2cd;
defparam memory_inst0.INIT_B = 256'hbbeddb94575b7ea8558f8b25f80c40f52bb92a098a0d87eb689710a88c0e34bd;
defparam memory_inst0.INIT_C = 256'hbdfb7e06c1918548bdaaf3904dceea50d7c73b55f71e0c069dbb40b47802a1b1;
defparam memory_inst0.INIT_D = 256'h20d3f5425aa39741f6285ead25cbc27e70388eada00b9cd68d1c9e4fb5660265;
defparam memory_inst0.INIT_E = 256'h82aa2c7d6722a7b4a3ce9c153469d028dc61889ac134cb1ac00c65c869ec2aa2;
defparam memory_inst0.INIT_F = 256'hb58658550faf454e77f0953e16568e846d5040a3896f5a1e30713416bba7c6ba;

Memory memory_inst1(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[1]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst1.INIT_0 = 256'h8d2a1283d7ded2a6d4e8dff6cdfe2ffdb798b76a284c4cd7bea325be2a753f69;
defparam memory_inst1.INIT_1 = 256'h193d622906e40f3807448e5706f592e1e2d525fd20b701ac000aafbc70c49e1e;
defparam memory_inst1.INIT_2 = 256'h82223d7dba4aa7bebc3631c2599fe6e8bbb37d3c1be13aa48125da6b52d9996d;
defparam memory_inst1.INIT_3 = 256'ha873f5b1d7597c9e33f17872bac18c0b863d03805353ffa25ca4d73f010a6404;
defparam memory_inst1.INIT_4 = 256'hcd82dddb6dcffcc4e12c8b5716b9e1e5b226033faab27bbaaaafca8cf69a2d56;
defparam memory_inst1.INIT_5 = 256'h61269c759f790a8779eac25af0634a951dee3b28554a1a2d3a3167a4914b9b44;
defparam memory_inst1.INIT_6 = 256'h93dea02bbd6fb74789c362aadf9d8d75501a765a343dfcd6323b99fb26f2c151;
defparam memory_inst1.INIT_7 = 256'h5393137b13f60695190a400b2d67e15f0b50599923c6ea2e494d2f84b4531cba;
defparam memory_inst1.INIT_8 = 256'h7d889adf0df0b04a50bdd3b17d35234cabc3287c9bcd7a9fd320e7d8edfe7393;
defparam memory_inst1.INIT_9 = 256'h5e8fcf125c218269ba471f44700c66215cbc84858c3abc1329df6c7e1f7f649d;
defparam memory_inst1.INIT_A = 256'h6ba6053287a49e5a074f7bae33167a198dc72a7afc37fa703ed162e3c516dde8;
defparam memory_inst1.INIT_B = 256'hfa3e43a045a7c04cc1225b17eec8db1a0755c21508c1da8d04349258fda59af0;
defparam memory_inst1.INIT_C = 256'h907daaf88f9a90584ea4f8c89152625868450cc37fb9a50ce346d4f84858472f;
defparam memory_inst1.INIT_D = 256'hb54eee3ccf3479c7d180e4bfa8f31966a40c1d73ee4107e8877d1375a2aa205d;
defparam memory_inst1.INIT_E = 256'h75207f5da11ef5e3da743ff932f0d367ff55e72c34fccb6119677253dd5a2844;
defparam memory_inst1.INIT_F = 256'h7747f311a5a45ee6baf56aeb0bc7535740029099fec36642d4f20b62ce6a3de0;

Memory memory_inst2(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[2]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst2.INIT_0 = 256'h57f9fd5f417f4737c318561fdaf4c3891fa780d601fe7bdd061dff1c11dca3ec;
defparam memory_inst2.INIT_1 = 256'hd12f20bacd7bb78745a66136e273cdee2efa4b3981bd3c3443ceb1616300f886;
defparam memory_inst2.INIT_2 = 256'hb9b002c66334651763d4f91fcdb7436f745d18abbc16e33db88543dd28a24549;
defparam memory_inst2.INIT_3 = 256'hba8dbee63cb3f983e6403b3dc79470258cd648b3c4de93060df79f8f8d7d3e6f;
defparam memory_inst2.INIT_4 = 256'hc8569548413896b64d61c64404edfe1e83a5ead1087d04e374029b469f0643ec;
defparam memory_inst2.INIT_5 = 256'h4dd2b6c3e512b39f96f02c4a8ff5f58cf70fa801a9621583e7260a89181593ae;
defparam memory_inst2.INIT_6 = 256'h4a5ebe5f8e0c3b44d856936a026e9047d0e9d6917fac1c33afc6e5abfb7443ac;
defparam memory_inst2.INIT_7 = 256'h0572a0705bde2ed2d56fb8811914ba8694c191536f0c06709e6ad92b9f47a6b7;
defparam memory_inst2.INIT_8 = 256'hfcfd1efd2f2ae3f80019c3d26af78d9501d7683f72ec359145e6558d6652d3e0;
defparam memory_inst2.INIT_9 = 256'h3a4ef11b27df8fbabd4f0d0020ca30eca2719f73e338d8d57b84ebb993d859ed;
defparam memory_inst2.INIT_A = 256'haea808593a5cb36e25abdd3084c3e1699266302909d2ae038b4a1d0f44ddbe36;
defparam memory_inst2.INIT_B = 256'h44146b92dee067d95c09c97f89fb61c00fd167fe56a0b9d8b5b4d9ea0dc7a790;
defparam memory_inst2.INIT_C = 256'h27eaa2cd7d66588c256a9deb61cc6f6e1b65dc2b453d79dd4e966e3faacd268d;
defparam memory_inst2.INIT_D = 256'h0cb6f65b8d325e1bd017654ea127542ef31fc43ce701b86379eb97d15df836d6;
defparam memory_inst2.INIT_E = 256'hb0245f68a5bb99e95fe2c84b4b78081daeb88217535782427fd9068bfbdb9174;
defparam memory_inst2.INIT_F = 256'h6bcc10640c984c777e1d7e54add5fd28b5115be6c17414428ed9493fa915d9a7;

Memory memory_inst3(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[3]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst3.INIT_0 = 256'h447ab672a9adbbaf36d57b95d665f103081ac75fc87d779bcbefcbf07b18db5d;
defparam memory_inst3.INIT_1 = 256'hc845a27daa9103971cfca6696dedbed2c47cb41f849e4c92b8ecf1649e5ef2ec;
defparam memory_inst3.INIT_2 = 256'h153c364e4aa0274a59c28c787f51a44ca0783fc4da1c99cb030a49302ccab5d2;
defparam memory_inst3.INIT_3 = 256'h5950304b57158443d46f22f447c5074a5a4e295ada23d65c60b44b24d5344de9;
defparam memory_inst3.INIT_4 = 256'h70f298e8f281d0e2d1bfe2abfe482de12b36f97ce521a2853603c026095d8066;
defparam memory_inst3.INIT_5 = 256'he4ac5c6fe7fcf8b3cda11a8a9231fad716e490ab8f87dfea97e3e9220b9e46a0;
defparam memory_inst3.INIT_6 = 256'h0ee825f23bf3b972f6c2840be9ffcca773a9828958fbc3e479a011e90bc8177f;
defparam memory_inst3.INIT_7 = 256'h562c6677eaf214b90d59be6d5a321284ae93977bdc7f9b2bbd4da274c779ba31;
defparam memory_inst3.INIT_8 = 256'hcd2c3dc29897ee3c6a9afe36ea12fdcee1c32e5e3967e05d27d6c21b06f2ecdf;
defparam memory_inst3.INIT_9 = 256'h21d24378c3876b017948098124c266d17dec0cf56f9b1bf447544fd99e74f7a1;
defparam memory_inst3.INIT_A = 256'hde84b0f345a8f486fb9b71535ab63e8fe404bba9eb9be7d54802433561994697;
defparam memory_inst3.INIT_B = 256'h97151be9712e0da46722c1ed035686fe72e6a900d07894e27ca3834460312eda;
defparam memory_inst3.INIT_C = 256'h4764663921f87a18735cd2d28b77ba5e1c25d19076b2d63b110467de56ae97ce;
defparam memory_inst3.INIT_D = 256'h01848c8827f53e0d41be108f9572984e72a5f44f4d7e5c9bb229aa2005c42112;
defparam memory_inst3.INIT_E = 256'h41d28c8ca14704cdb15be2729cd7691de74a9ba2936d5a05a197c14a0717f215;
defparam memory_inst3.INIT_F = 256'h139433b5216d12620ccaa262df1c92286a6e1ead7d513c5dbb13aa0db342df30;

Memory memory_inst4(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[4]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst4.INIT_0 = 256'h51d5396a2ca53bfc87dc128763fb8885385d95b2c9d9c3711cf19738212c9e21;
defparam memory_inst4.INIT_1 = 256'hc7c97aa57175d868d0d9a3858f9ede4ca59316f3da92054c3d3599a79150c1c9;
defparam memory_inst4.INIT_2 = 256'h1861d9cef72a616f68a35c3f5a87aa00ee07b45624b16fbc12cc003e259c399e;
defparam memory_inst4.INIT_3 = 256'ha60be2de71b7c9dc9583b93e948a593282e9b45fd542b8405bb5c08cff79af40;
defparam memory_inst4.INIT_4 = 256'h05de1253cd9776fa5e3fc2a8a9fe72a833905ce5dd3eca7b2a29054de370a047;
defparam memory_inst4.INIT_5 = 256'hfe8d492b33289c1729724b619d653cefa5f7d599f2aab601b9ad67d19a043a6e;
defparam memory_inst4.INIT_6 = 256'h4087659c48cce1947e678942e005b1c0783882e4cc2db4b5cc38d869fbefb9d4;
defparam memory_inst4.INIT_7 = 256'he8bacf4998c4f5f1dfb665084fe1305cb14fbdd01c3a642ccadcd1d8b22afc34;
defparam memory_inst4.INIT_8 = 256'h9decc25f7c6dafdcf33736fdbde1b4274bdd6a948f16437d8bc7ac960e931958;
defparam memory_inst4.INIT_9 = 256'h06c7d68b3787f4687decc105da558e961025eeac4aabdf68ce3422166b2dcc49;
defparam memory_inst4.INIT_A = 256'h242d88cd4f42a10c23f511dee0be45ecc7f5d2c6a2da9964915c8de29130c53f;
defparam memory_inst4.INIT_B = 256'ha3456d1c03ac6e53adeddc9df55af72ffd9d3b1df960ff68172ce588e3f76b8d;
defparam memory_inst4.INIT_C = 256'h949e9cadf3852c6b04a3a465451f7a24a07cccdf650e0ae6060e1fa23b3f61a4;
defparam memory_inst4.INIT_D = 256'hac0ece782f9c256dbf76b8e9f54f35baeab9a3d3394eb17d2c6b490e3def47fa;
defparam memory_inst4.INIT_E = 256'hf660f29ea11bf431a239da1a61a11b65a6d871c2febf527b54d9b974a1b9059a;
defparam memory_inst4.INIT_F = 256'ha3c1bb72945bc3504c7db3d0d197295f935d078e0cee4a0fa432a453a2b6b336;

Memory memory_inst5(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[5]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst5.INIT_0 = 256'h14af041d02db615f84737b0b9a3001377d6980fada219a50e208d11117bf1d34;
defparam memory_inst5.INIT_1 = 256'h31ed100d46f5847e246a16f71cc41accf13eaa577a8157d22659539809ccfcc8;
defparam memory_inst5.INIT_2 = 256'h6179c9b479c9d0b6045d92207b9070576b0a3cc1712c321dcf45d05d6ba487c3;
defparam memory_inst5.INIT_3 = 256'hf5ddb03afe298fcb2d639ffddd88180a3f79d7bbffeca24b267bd086a8ed0c3e;
defparam memory_inst5.INIT_4 = 256'h584719ac49f7fefe02ab059ee39e3e27eba905eb311cdc4c82da4f05b7451a9f;
defparam memory_inst5.INIT_5 = 256'hb7eaa09e05efc0e08aa0de024aed17c1cd90e8a548c1e86880e8a00bce53e59a;
defparam memory_inst5.INIT_6 = 256'h6fa017ec1c8d711e22010cc634069904ecbd0fe43bf97482db0301b0b24f38bc;
defparam memory_inst5.INIT_7 = 256'he27fcceddb7acaa5f6f9c0bda4c14f305231aa227a447e49d4076331f9f82ac2;
defparam memory_inst5.INIT_8 = 256'he16e9dab740c64a39de858312216169e362e3c99eab0870f3c04a58cf5c5d822;
defparam memory_inst5.INIT_9 = 256'hb1978cf97c50fa3b64f1bb46c73e5a4eece7217309211847ba4dc711ba335bf0;
defparam memory_inst5.INIT_A = 256'h407ebba7fdbd3154e2e3783e5cf5960396e5dd854709476da7871c428f3d9c8c;
defparam memory_inst5.INIT_B = 256'h747609f17238130afc02edcfe15f7c5d5f8a7859d841b119406ec0cdc7c0a61b;
defparam memory_inst5.INIT_C = 256'hc8f0aad680ef6c9e0a3c9965ade9e7f13c51cd70369ac00edb2405e06210549e;
defparam memory_inst5.INIT_D = 256'h58da32bd6659a05c3d2fcfb4a4d193d5fce175d6ea66b0a5dc0d4a54e7059db4;
defparam memory_inst5.INIT_E = 256'hf2bf1d18b6ace9d3979eb1e2cab53c488e81853d3054d0cc8a89878e3a0ccd7d;
defparam memory_inst5.INIT_F = 256'h762889929f13d6946ca9ab9653ac84d9ce30c4ec273a4e2fd5e1642e3eae5a4f;

Memory memory_inst6(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[6]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst6.INIT_0 = 256'hb36f3f74256503fe2980edf8a7908e1b491ae7797f188b90b944be086e8e95ea;
defparam memory_inst6.INIT_1 = 256'hd3f21b7146a5410aa0d3c2474a51823deac5a906ab03af9ab7b61d84e2ab5c7d;
defparam memory_inst6.INIT_2 = 256'h9747d3407041530ee9c871e5b4d7ff94618d85c62341781974f6226c3841b9f3;
defparam memory_inst6.INIT_3 = 256'ha10c3360ab434d4b719412dfd9dbd4474ca3b167c254dd212d45d8c195ff8400;
defparam memory_inst6.INIT_4 = 256'hb52d61df47f571125993b8ff7bed4be5e7fb4f853135bc22c71f2040c33a140e;
defparam memory_inst6.INIT_5 = 256'hcf3dab94c62732c7662b3593a79809b59bf4c75c4cfd82b0df64af7f47437c7d;
defparam memory_inst6.INIT_6 = 256'h3e3ef7355e2f189963200cf49335b50fea28c33862683944cad8644eb47b9b5c;
defparam memory_inst6.INIT_7 = 256'hb9b1a16a54edad1cb80deb7a95563525511b9221983d8884ac26257761d4fd85;
defparam memory_inst6.INIT_8 = 256'hac1efb59ad1217048b730209bc458136cdefce76ed1d75694b6bc400815b4a1a;
defparam memory_inst6.INIT_9 = 256'hb49f8e9661836e450e137a223612a7e70ea040f73b36335dc3ddd5ad296425ab;
defparam memory_inst6.INIT_A = 256'h27fd86ce99a89177d5c36a65e98cde7e1a0aabf26fd22299021687d7f313611d;
defparam memory_inst6.INIT_B = 256'h1b120ff0c3868124f5d3ffe3447089770ed221a45dae24096573f1eb468d655e;
defparam memory_inst6.INIT_C = 256'hdc016bc017e48118145fd6b6ae18f0876f1c7b4f78c2048593798d601b05df71;
defparam memory_inst6.INIT_D = 256'hd636045cf77217888778ad32ac8c2429886e4cfe6fd294f82eda1cde4ec71b0b;
defparam memory_inst6.INIT_E = 256'hc2b938e43d9aa0b3843e61466e14fdc28684bc7539fd2dfac0df172951c344b8;
defparam memory_inst6.INIT_F = 256'hcaa3fa500a77165953388fed36039babd12bb93f13f45558db36dfbab423cf08;

Memory memory_inst7(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[7]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst7.INIT_0 = 256'he0c33d37ad8580f4ab56b176f1e43c3e316ded508e76681db2ec07d1dc393c3b;
defparam memory_inst7.INIT_1 = 256'h96e754111b6da59558bf16828e88b8e1dda3c69a6cd319b1010235d1bc3e3737;
defparam memory_inst7.INIT_2 = 256'h54280bca96d59bac2018fb286c8ed1176c6c4615d04bf992ed728346f0858bdd;
defparam memory_inst7.INIT_3 = 256'h60988e9f13970c3968263431f3bf76503cee6839a60c00c13e4d33f2f4c7c80a;
defparam memory_inst7.INIT_4 = 256'hdd49f19c092884ed2e03169e7ac503d154e11d9631f19de9c1f35553198c8939;
defparam memory_inst7.INIT_5 = 256'h59e59369516114bcfa80f9cf6151f162e405109ebe49e40204154d898309110f;
defparam memory_inst7.INIT_6 = 256'h74a71ff969509bda3bd5f7e45f4ea8212cdf141af488c71f18a75d517003cf8c;
defparam memory_inst7.INIT_7 = 256'h667918174cf10124eaff5728b69099e782a6933bff042b9e8f7fdd4096630ab0;
defparam memory_inst7.INIT_8 = 256'h8661004b3aedde719d88861d72e6985f1282d3a8f746189c1951b7f1981d7a7a;
defparam memory_inst7.INIT_9 = 256'hd71ffafc0134957643411554595a0bf79a91917523ef9a79c7639e39c8c4be57;
defparam memory_inst7.INIT_A = 256'h082a608e8192499a2bd8b8011095383d14c80e4143d7f521530a132ae4cbca90;
defparam memory_inst7.INIT_B = 256'h73c532f38711876b638cc0f2c24da1d88b9f639a8a16450e980ddd1fe923af13;
defparam memory_inst7.INIT_C = 256'h050bc97a5ee86c19c4e83fca317ac879d0ed0b919fb3a72bdc384c7302a56ad8;
defparam memory_inst7.INIT_D = 256'h378f8ef827bf40e7b2cd3b479d74d12202eee317ad1c3dc943efe7298eeb2c14;
defparam memory_inst7.INIT_E = 256'hefff49f85f9d83c1e4f7a4683d7e6c64b31ccfcf812da4b9a0ad5947025d8e6a;
defparam memory_inst7.INIT_F = 256'h00b1cfca9db546d42d78b3d107a9219671ce0d0ea92b819d3c98deb35fb09b62;

Memory memory_inst8(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[8]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst8.INIT_0 = 256'hc64c7246a0e72af1f4e7c81d2f3f637bbd0f9deaeb1e17d4f4e2539d2d6220ea;
defparam memory_inst8.INIT_1 = 256'h9492d547570c44978ecb27cd2540d4a3bf99310bd8de384a3afd5a370da977d0;
defparam memory_inst8.INIT_2 = 256'hbd4f31707ab1c7b5d226f9a146e60d226f0355fdff6896cc20cda208762e44e5;
defparam memory_inst8.INIT_3 = 256'h4c962f952335c8e3bfd9c2632c406cf2923979e5e3c30c8adcf028eb19d0fb62;
defparam memory_inst8.INIT_4 = 256'h7ad7782213fb02ac931fbd076187ab88c98eaa7323a861198e68d3cf59e919ba;
defparam memory_inst8.INIT_5 = 256'h6119cf7f9d7d10305701cc1c982dd69073cce44fc674a5e871dbd08bc1366b9c;
defparam memory_inst8.INIT_6 = 256'h01b5e1a61d90603c9ecef572cdab649fa8d91b957829f9efbc9aa9305b9dad12;
defparam memory_inst8.INIT_7 = 256'ha75ab41ca27e7b4640561c174d0de6a81837644c183f0d9366dd03e28023c0e0;
defparam memory_inst8.INIT_8 = 256'h5318509fd13f0eac05289ba81c0a7675b4f1af49ac70ebbffb90cc5ebb2fa053;
defparam memory_inst8.INIT_9 = 256'h1950fec04f595b52b4397808e6ce15c339dbc0de70bbe58999ac736f9a91c942;
defparam memory_inst8.INIT_A = 256'h346945934f003796d3b8c5432e8b823b97670be7c02139c8391439d154b5bb62;
defparam memory_inst8.INIT_B = 256'hfd088554a2aea2ac3917210b5442456c4d37470f43d445cdfb794ca39dc70eac;
defparam memory_inst8.INIT_C = 256'h38143763e2f88230268d5b2eee35ff707eecd68eceacaadb39db79cda2368b9a;
defparam memory_inst8.INIT_D = 256'ha9a4e21ea5ef67f7d44c976bf07fc6cbf7a35856a93499f14082beaf47c03813;
defparam memory_inst8.INIT_E = 256'hc18d42d3a1b1c662dd6d480b6835509c08a2c5a8d1c2edd9fb7d6529f913fbe5;
defparam memory_inst8.INIT_F = 256'h04cbddb6df87fed8b817c520b299b6e826454adbc6f2e5d853c53f9abb5cfafb;

Memory memory_inst9(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[9]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst9.INIT_0 = 256'h9c605f1a492ee25e28ef5c78965bf6a29a4e8d401cc3a83a2fbe7d2db9791faf;
defparam memory_inst9.INIT_1 = 256'h8126c922bb01d32afb25706b6f839969e9a9954cbb087790f92e9135f079d387;
defparam memory_inst9.INIT_2 = 256'h113d73396cc53214b7757c36890c7493d828c2417fc632c1faa688dd134ecbfc;
defparam memory_inst9.INIT_3 = 256'h46c8b3f111793edddbcf8da43668510182ec833e84ddf79f3a58c0cfc800b555;
defparam memory_inst9.INIT_4 = 256'hc0a371c443dbe3a187d3c98abdcec22054bfc818b86b9b21818e343e23792957;
defparam memory_inst9.INIT_5 = 256'h6974678354a639151a9baef7cf0e9efec7c650078be6dbfcb677798206dfcc16;
defparam memory_inst9.INIT_6 = 256'h65cbf766018783d22d46f70b974efc0aa3f27e9db3951d1a037046cfcaff5928;
defparam memory_inst9.INIT_7 = 256'h55b6dd55e433f97b67cc949f3e32fac1aa23e60ae713892f9db94e8bf917e25d;
defparam memory_inst9.INIT_8 = 256'h9e6a21de9f572ee48ed8832d8006aef048cede81b2f76d337d4bfac6b0d60e3e;
defparam memory_inst9.INIT_9 = 256'hbd776045653d89501e5206e50a1de888c2d3733c117b619c2d6eb1a4a952a2b0;
defparam memory_inst9.INIT_A = 256'hf1b11e495b5335a7cbc5f629b4f4f3df6dc6c7e4b2604d59d8611c132c2c3a6e;
defparam memory_inst9.INIT_B = 256'hb9283849cb6dd1f3e43fd0979fc6044c0dd8e3a24b95a0a16a2fea8d255aaa1c;
defparam memory_inst9.INIT_C = 256'hc987c12fff169cad086d5489faa506699f9a169c73fd55ac1dd21d0a84de6d99;
defparam memory_inst9.INIT_D = 256'hb1761fcec729b1c8a18d6a35d8fffe6e42d32ab4ab049e3f187af1c9540de74b;
defparam memory_inst9.INIT_E = 256'he463fe056e86075804b1c8d186655ee42c1c7036c278bce77ee0946d77d5f0c8;
defparam memory_inst9.INIT_F = 256'h92b8a17ca8232b523e4249af35fa5bddf015b4b2909906d048b3c5a574318e3a;

Memory memory_inst10(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[10]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst10.INIT_0 = 256'h7f72915a6c007ddf14ae86d192c61b50bd621f5e417af588684e9165c894d83c;
defparam memory_inst10.INIT_1 = 256'h082a275dd28ed6f9448045f336f0ee3bcf205a3b5a0a4c05477b548d00e16e09;
defparam memory_inst10.INIT_2 = 256'hdbc73b0afa83ef2f2c0e0fe4eaa49e049f2d5ba5439932e81f13deafaa39716e;
defparam memory_inst10.INIT_3 = 256'h3e5c4591c1622eb2fea7682ed3a934fadb6d0417e8b0eb0199e6bb3af8ae0e20;
defparam memory_inst10.INIT_4 = 256'hc7a2c22cacf7f460fd785bc7dbe78be33becdfb76a77adad19dcbbf28903cf4e;
defparam memory_inst10.INIT_5 = 256'h8fe96fabf08bb1e7b8be390ae531126b518601390fae2dcfa49e07839a3883fd;
defparam memory_inst10.INIT_6 = 256'h1dd242dcb0e24fcbfa87fc9aae24af3380f147774f4574247fbd64d918ca4a3a;
defparam memory_inst10.INIT_7 = 256'hea832544cf516ca131ed5f34c0d81cb82d2b84b6329904a22e8b5ca6ea362ee2;
defparam memory_inst10.INIT_8 = 256'h85f81abd1d638a13a69b1096346bc69539a17e55e0a5a765379c36301bb5973d;
defparam memory_inst10.INIT_9 = 256'hb071bd091ece0a1b0ecd62505f9cbb3819f511d99a1d5e955716544a93ca8457;
defparam memory_inst10.INIT_A = 256'hd7ae78db43fd39ebf917814e5513d2f768f2b86c53c2e0322692de2286fddc26;
defparam memory_inst10.INIT_B = 256'hc28681ba425959951a983c07658690647b733b635b403b2c81f1286167e6fa50;
defparam memory_inst10.INIT_C = 256'h370dc4d2371b6421927b6fcbae8e1cfb82d9caaa557b657c5ecdb88609518604;
defparam memory_inst10.INIT_D = 256'h060707d26aa9c6f0bd6e4d1af2a9ebb79256a22d01d4bed5fcab4e70099432c3;
defparam memory_inst10.INIT_E = 256'hf6f5bb7c55890db61759ba64a9f2258b8beade693a13c7ff37d311e851cc43ee;
defparam memory_inst10.INIT_F = 256'h13b744949beb787de859ded4a16858560c536f84ea2387c353fc5cc88ec6e132;

Memory memory_inst11(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[11]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst11.INIT_0 = 256'h97028312bf212cc03dba20a26daf7918ef377f6211eb7ed67ed829a170d8622b;
defparam memory_inst11.INIT_1 = 256'h55051ea504b3aa821bbc96e791c6e4d3a7a0d4d288ad53b1a84b54ac941952fd;
defparam memory_inst11.INIT_2 = 256'hfe3a6f1f5b28fa838d0cf0315dfdb0e2df9a7a67e4aaa90135f463c9e525a60c;
defparam memory_inst11.INIT_3 = 256'h7768758ed46ee3a3826f6fd4cdcdbf0d4bca58741eb1f6e376afec05f2ff910a;
defparam memory_inst11.INIT_4 = 256'hc6eeb079024212549da225693107830ec9ded4cde7113e5c052b914f42c13482;
defparam memory_inst11.INIT_5 = 256'h3fcd05e7ed13510b14960c0aec73e832ab7a599c2e3f6c8e63c51600dd9857fc;
defparam memory_inst11.INIT_6 = 256'h0cb9e820a73b758be535ef4a0ed796eb861c67fb94a7786997c400cce022ab76;
defparam memory_inst11.INIT_7 = 256'h92d0087adc97daf77c74ba36a7316d5459ff622fd6c14aa41fb909382a7eea24;
defparam memory_inst11.INIT_8 = 256'h4bc38670d43263c8e1164a555351fcefb9caf62499ece08b5250515edc665b49;
defparam memory_inst11.INIT_9 = 256'h513299739757b4b510c3043a425588422f87519029654c2754fb59d9a40df53a;
defparam memory_inst11.INIT_A = 256'h2f301b3394ec4156ee45ee4b30e2076fb715a228c5035eed35ec7595de340d4c;
defparam memory_inst11.INIT_B = 256'h67b56c945b4b41da55eadb2cd4b3f21bdec4b9b06212efffdf157135d6432faa;
defparam memory_inst11.INIT_C = 256'haea6728e301b55c9b8fec37c0d5d859e92f165c595cd5d4143219f59bcfa3542;
defparam memory_inst11.INIT_D = 256'he887e7f90e6d9dec47fb605adb0bf32331c327b0f4202cccdcf83476a6272ce8;
defparam memory_inst11.INIT_E = 256'h76fa65bd7152ce719f30d6178e5d8262d0c3e80dba778db35da442dbd235b11a;
defparam memory_inst11.INIT_F = 256'hee048f75a0e8f97a9463213adcc62d5358ca021956d0467d423429f371ee36e4;

Memory memory_inst12(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[12]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst12.INIT_0 = 256'hbfbbc7cc3ff62d3a769223e5c1edaa86d3e6e8a5a62c57a5bcd3380288885474;
defparam memory_inst12.INIT_1 = 256'h24c153275ef11bb77f4288af1ab2f53df27617cb231cb7ab83bf3fd1a3cb7b82;
defparam memory_inst12.INIT_2 = 256'hc6b3209465fbe7218894249962cff58eea6f452e42a7574f645a8de94ae03961;
defparam memory_inst12.INIT_3 = 256'h9192cb66e81c1281c694e1bfcaea713a82608dbf89164d32718cd823b386d968;
defparam memory_inst12.INIT_4 = 256'hfef0dd6f016d0859795d2a185d8be41cdc9bfac32fa9b6e42a3f32417be63bca;
defparam memory_inst12.INIT_5 = 256'ha7e957c495a02afd8ea228bc4c168d5f2210e0655a20a928d64026f0498e1521;
defparam memory_inst12.INIT_6 = 256'h4dc2b208977f5ad41309b24fb349d316c2e12bdd0fcca3598dacc17fc043546a;
defparam memory_inst12.INIT_7 = 256'haca79b086f9602453fb5dbef27855b5ed1f9d117c39557807d7e29f7fce5897b;
defparam memory_inst12.INIT_8 = 256'hbf2b911dd336638a4fa93f03acabb94984425b72b9ff2e617d8df28f4e8240c0;
defparam memory_inst12.INIT_9 = 256'heaa99fdf1bb71a34b11147b6728bd804ac58041cdfe71ad338ba04c0a91cb6e3;
defparam memory_inst12.INIT_A = 256'h0eb63d5891074c844c7eb0251296c168080123fcf5d72548b4282483bef5072e;
defparam memory_inst12.INIT_B = 256'h250d0aa79af9a81a62075a3dc72b96a44abb266818eb2bfda9c0f6757ec5598c;
defparam memory_inst12.INIT_C = 256'hc6b9ea45b16405d7b0a6ebfbe37c98460a40226a55c8a53bad062209cb7d237f;
defparam memory_inst12.INIT_D = 256'hed40d10df0e8e0bc71389bbc2e1e2c13bb0315770a0d121aa28ef0a3c199d6cc;
defparam memory_inst12.INIT_E = 256'hab241fd1222be07bc241bd16c42465e14944a5462ef16e794c8035f8f0706ed0;
defparam memory_inst12.INIT_F = 256'ha199cdcfeefdf0ad9c09e568a995fa44c38fa841ebe28f81467f6fae1f4bc19c;

Memory memory_inst13(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[13]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst13.INIT_0 = 256'h01a71213be6161df14c5f964b4a92e1b4c55252f2200baa57094af96d66f6c19;
defparam memory_inst13.INIT_1 = 256'h893a5abf59708d8b930c39703377a49fd572c4abe977ceea660b006fea9c3a4d;
defparam memory_inst13.INIT_2 = 256'hd1ab277864b04258cd6fea484e1958d4410df3bb80a9c06d7961b43213232557;
defparam memory_inst13.INIT_3 = 256'he777d0c8c034c59b429e7bbb7e169b7cc7b37ada63155f4bee18d6e54f9f7410;
defparam memory_inst13.INIT_4 = 256'hce3572f8cf57b791280aab771eaa005a80aef51ec803c0110f4bd40a3a7e2e26;
defparam memory_inst13.INIT_5 = 256'hb17da02cd4eb7ce8e73be9e14c1f9e9bcd27feeb6e283848960a39da59db0ff9;
defparam memory_inst13.INIT_6 = 256'h8bb36a7fd61acae1f4e021ef6cafc526755c5d3735cbabd2f1cfbc7b0c5124f7;
defparam memory_inst13.INIT_7 = 256'h064ed4b939fd0f156b13eb7ce2adc39c95d2709187b643843ed27e3244cb2ce5;
defparam memory_inst13.INIT_8 = 256'h988826caa716ceecf610972d7ffdb918347d2cee3d18fd9e81bb91f85789fc95;
defparam memory_inst13.INIT_9 = 256'he1fa180363067a6a37a730fc68adef17e700b4c257324c0df3fbdc78f18e4bda;
defparam memory_inst13.INIT_A = 256'h7eceae8888247bd450b6c8c66c21591420d20d2990915a951d5b1b4f79820292;
defparam memory_inst13.INIT_B = 256'h000ea0fbd6e603baa56a58f5c1c83065a7cf227c58e96b3ea84d71a15f434831;
defparam memory_inst13.INIT_C = 256'h9cd9f692b9aee976df614fb29bf0a797eebd2c67e5193a9ef7d75bfb3db1635d;
defparam memory_inst13.INIT_D = 256'he549c27d803b36095c3b8bbb531a7b5b8fb7d9f8c9542f7490338487b461a9f7;
defparam memory_inst13.INIT_E = 256'hb3e3f299a831cec89d7bafda8d979f278c2705f06cd199efb9bb7d3d0910264f;
defparam memory_inst13.INIT_F = 256'he0e3f352e6c71852ec272b43916abc0d1cc53cb02ef29b515d27d82739d3c71c;

Memory memory_inst14(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[14]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst14.INIT_0 = 256'h87fd56ea9f1aaed39f57b9b47a8b30513692a1c86f234e03f127723f35a42b81;
defparam memory_inst14.INIT_1 = 256'h27e12683a771a2f7b8d987d71203e1c72c12042332dd9ac9c96015e7559cf13c;
defparam memory_inst14.INIT_2 = 256'hd5fff20fa48c77675bad180ed218e63cc89e65fbfac53231e5b8827d92f9b655;
defparam memory_inst14.INIT_3 = 256'h64c27c45c443c6b4c429d7b501742de95d20a0ae209d6bbc146b87341fda5dd2;
defparam memory_inst14.INIT_4 = 256'h62348aa0ce5412423673f6b0a0b9adc608c76870cf3b4ca865b328c67f685c17;
defparam memory_inst14.INIT_5 = 256'h9d41c2fc2ac5bca4e0890286503f823e843d54812c77335c8fddc1aac074a479;
defparam memory_inst14.INIT_6 = 256'h58584df4b72b1bdee4568cb3391af284e94f7ea981514553e88bbc4420d41202;
defparam memory_inst14.INIT_7 = 256'h72aa593239dd70f9bf2f6162874473adb2bd093fdeae25d5abd8be9b885596bb;
defparam memory_inst14.INIT_8 = 256'h84bda277a06a235c2b120e827e3ac296a50ea1e3c79662662627caaddc09403d;
defparam memory_inst14.INIT_9 = 256'h478a55f6b8bba47113ec49c314dfe5fc72d12dd5008202204b8e9f2e5606d2a6;
defparam memory_inst14.INIT_A = 256'haa7624700064a7b176c02de8d49da65a31d3844b766052c6c8fa873b55374f18;
defparam memory_inst14.INIT_B = 256'h950a1317147b46c2802220b32cf5c60e505b09130993f65383b7961f1848a4d0;
defparam memory_inst14.INIT_C = 256'hdb4f98ff405ffadc503c88f4bf6489f4bcc9095f21026b2cadb631ec8aa37dc6;
defparam memory_inst14.INIT_D = 256'haf43a552263f5a8301d86e8edd6fbfc34b830c65ed840ade3d595e21db90deb6;
defparam memory_inst14.INIT_E = 256'h97ab84509d2362b4d1305727a268da8c6fa44199b1bd1a377ef068acbb5ca3b7;
defparam memory_inst14.INIT_F = 256'heff1b3700bbb7b40b29ae77f85d4cb67592e58699117f45fdd2ecd746c90348d;

Memory memory_inst15(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[15]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst15.INIT_0 = 256'hd38b4b4aa3ba90d05b9dcf58aa687fb88cab44006dde84712862a0fe5b384e87;
defparam memory_inst15.INIT_1 = 256'h30c6c86dc71c3c384a5d7ea8b7cb502b4547250c26bf302a6272c1550fe0c71d;
defparam memory_inst15.INIT_2 = 256'h26d5922f4919b392f45e9a9628ed94034e5f75b3b6ac624a19e55669c320b47a;
defparam memory_inst15.INIT_3 = 256'h4c84a49cb61f3355ff70dcfd1fc96d7aa2bf468512e5c3de8a759d8273a21bab;
defparam memory_inst15.INIT_4 = 256'h95f55509d76369a00074122dfa3b527dfdcf43075608eb2588437f46ea17f69a;
defparam memory_inst15.INIT_5 = 256'h1d6d925aefd9e1881807732d5bccbb009265dfc0afd53b97f3fcfff9da52877d;
defparam memory_inst15.INIT_6 = 256'h77585b7dcbee17a3f5e20dc1e4d5740e651f8b503447e5de62c642817c172b52;
defparam memory_inst15.INIT_7 = 256'had003a0e9ff29ab41466f3ec7c575afe724a909f27e9d9932e411f0a973344ea;
defparam memory_inst15.INIT_8 = 256'he39ce0a39e6e3163ed254aa4300429f0f9265016614298709b4b166467b1921e;
defparam memory_inst15.INIT_9 = 256'h5af43b537bd2338c1bd0752da7916ab10d95ed7e91f75b6fb29fdf100ef8b5de;
defparam memory_inst15.INIT_A = 256'h1ae2bb3754d3f316597648132492d8eb5a8871ea32594cee4be4b416bcedc03d;
defparam memory_inst15.INIT_B = 256'h7de3d80546b4775ca5f21515fe2348dd7b4389166993730bd6241e3f3230445e;
defparam memory_inst15.INIT_C = 256'h85145a918395627867082e02f7f51c4763a653b3393d84e685ed06b5a3bbef9d;
defparam memory_inst15.INIT_D = 256'hd58027a637cf4d41d0eb63a5d0080751bf522529165b18cec16ba721d13ea34b;
defparam memory_inst15.INIT_E = 256'h36cd39c5f6f3669c30fbb368d98d80a695e39b697f1aacc147ec0b2394a1cdb0;
defparam memory_inst15.INIT_F = 256'h9aca4927e89196c00a6ebe99997a8d94d7f8578e3676cf3839868c9934afff5c;

Memory memory_inst16(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[16]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst16.INIT_0 = 256'h39e2d2fb929f6634fb850ffcca5380a1c2ba7644c664ac57413a2fb2a89a81a3;
defparam memory_inst16.INIT_1 = 256'hc19dbedceddc24f37fd1171f68b8cb949c63215f447e83a55befa57c54256dc4;
defparam memory_inst16.INIT_2 = 256'h56c584664d8c2a6e1b7294ad291ae51890d75a18a84ddb0ef018bf54ce475aa1;
defparam memory_inst16.INIT_3 = 256'h578f8d76b8db58fe026bc36e80e1dc455f2636b28559191ca441c84b8a5e7b09;
defparam memory_inst16.INIT_4 = 256'h9acd5f9b72375915182c462b5525230bca77ec57ef991ae3bd576b9ded55611a;
defparam memory_inst16.INIT_5 = 256'hea082a5c36e2959ae05fefc9d1d59bf966195738eea111d226ee413352ca3503;
defparam memory_inst16.INIT_6 = 256'h934d8b34b76fb090a972c3fee8e7f00c51941f7e449ddd94fc3bd2d11c940809;
defparam memory_inst16.INIT_7 = 256'h4eb87167e908e5c42b3a8ada1f95e700c3aa691177df240e686e1499398d7345;
defparam memory_inst16.INIT_8 = 256'h9234ab5f3ef2d26da0db963e895fd774591e72c5a571b43a520808b01e9ce930;
defparam memory_inst16.INIT_9 = 256'ha6ac0fd5b0e51646ab158f776511e760d3175f702622b00372c4da899da3c882;
defparam memory_inst16.INIT_A = 256'h2f7d53ff83e71ad13a0e562abaeffd6b5711cebf12e506de52bf7859cda180bd;
defparam memory_inst16.INIT_B = 256'h239d3a3cbf06ee442445bd05583ece8f8b8f1042840ca771c05da9e98f848707;
defparam memory_inst16.INIT_C = 256'h7c770c08f730946456c805b039e7c606ce804051f896168d454f1f69d3a43f4b;
defparam memory_inst16.INIT_D = 256'hc3ca8910335f175db56d0479b157ea1b5fd2f4646a831d94d6eb811dc6195112;
defparam memory_inst16.INIT_E = 256'h97e3e1c1f0b6483fb5e9a9529e0cc70072f24b12ad9c6c35bef77c11ef0c7afd;
defparam memory_inst16.INIT_F = 256'he45747933c426126382ebc62642236a14dbf3bbf33b10ef323e66af58768442b;

Memory memory_inst17(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[17]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst17.INIT_0 = 256'h5bce46d4fa0fc575b92c77085a9c93783a1b6c5e943171d02792cea24652c1f2;
defparam memory_inst17.INIT_1 = 256'h4e9addfcbfbbcf05aca7c24f307bea9d443d950727249c65ffe800b826fd8059;
defparam memory_inst17.INIT_2 = 256'hd5519f3f79851a50a979ff8bccc73abf62fed27dd31fadea7a84261cf2870a43;
defparam memory_inst17.INIT_3 = 256'hb98a230f9db9b840d5d510592b369af11bdb5d4f4d0fbfed20a8eda00a7582ed;
defparam memory_inst17.INIT_4 = 256'hce0f5a6a6b29af90fc26fd3db766dbecd28cfc2cd865951ff9d31b5a38217d9a;
defparam memory_inst17.INIT_5 = 256'h41e9e018a5eac6bee4b59cde2087e8a907802708955369c54906cdd5242260f2;
defparam memory_inst17.INIT_6 = 256'hbadd060030ca5bd04e3e4678a93c11a16b63fa02e2c2017fbeec46bb7d7a9087;
defparam memory_inst17.INIT_7 = 256'h938ae4bd03b401a8b612a3af7942d8ff31fc2d09ed0f32e28577e2a916fdd33f;
defparam memory_inst17.INIT_8 = 256'hf581d12b60cd1c5f25a76c74a9a2d9405ddd2b20f8330f4faf660fd71b45ea33;
defparam memory_inst17.INIT_9 = 256'hacd707871dce7418fb1551483c710a8e41017f4d43e6b55fc5c90900a09b713c;
defparam memory_inst17.INIT_A = 256'hf63c49cb9574fb5cef381c713390d6d47d4ddf962b240888e66d401ae0368b58;
defparam memory_inst17.INIT_B = 256'ha0968ad5193079c85974fcc26036d3fc169d56ee66dfdb34bb88559e9930f388;
defparam memory_inst17.INIT_C = 256'hd5829dac9f3cab4774d792fae8e3188afdc07f73cd71d6999c068de19b139ca2;
defparam memory_inst17.INIT_D = 256'hcdbc994f1b3a942acebc6d3180e149fb78c919e612ff04a112cf4c37e718fc6f;
defparam memory_inst17.INIT_E = 256'h437dc7f8a34a633815c481e73d2fc2fdc3b0619b9830d23eadc74658516a1468;
defparam memory_inst17.INIT_F = 256'h9d9cbf8939c9e3f767ed07cab3397f0777e50eb4219532cffb404fb4ee22ac2a;

Memory memory_inst18(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[18]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst18.INIT_0 = 256'hd9e14a50eb06758eaef7d024fa59853c42505fdf045d78208bf898e1466a19ac;
defparam memory_inst18.INIT_1 = 256'h83f2886951841dfd3277c17aca6a187b34ff78ee548d8801d4d5e625d46410f1;
defparam memory_inst18.INIT_2 = 256'h94e366958f44d640d4bf739de3b9f868878703de146709b14fd5c0f57fea37d7;
defparam memory_inst18.INIT_3 = 256'h5c4fbe36aa7615092a03dfa73505c12aa6da90b5b0d4fa7c18ef08fbc931bc58;
defparam memory_inst18.INIT_4 = 256'he522364ce9ded1f27d9d846d9896d67c3ff8cd6b02b15543fcd3771b0aeb645e;
defparam memory_inst18.INIT_5 = 256'h034f4445f2635c6c8c9e2cd126befcb0ee17da695b7ff52137d461dbf6bfadf0;
defparam memory_inst18.INIT_6 = 256'hbd8d60ffbd85a00a40a6ee7fd99bf4d412425247cd0ac522f1b55d57c91c97d9;
defparam memory_inst18.INIT_7 = 256'h3bff463d6b54b68be2c561f0ad83547c291f4ff0e1301d43976d077f95938682;
defparam memory_inst18.INIT_8 = 256'h9a0d96ad60bc115d1a63bc1c2c96db587f5a8520eac99f9c98ace03a26fb6bbb;
defparam memory_inst18.INIT_9 = 256'hbb01a3911e769cdcf291c3b1c5398addfeb18ddb33ad624bc5a682875ae90549;
defparam memory_inst18.INIT_A = 256'h6d35db9a174701000e56bac90c4cf71a210d015722bce06fe1f6d7ab417c2728;
defparam memory_inst18.INIT_B = 256'hefc4f06a323c3e843d0d61101f5ac2ee99ccb6b9c1806518e88a60220197484e;
defparam memory_inst18.INIT_C = 256'h3ada433c4a7a85069db434dc4526ad4133227adff96b3fc8b4d90e1accd7668c;
defparam memory_inst18.INIT_D = 256'h66e41ce45ceff73c70f962d02abe06749f3b779a89f8b3894205ab40b41ee4cd;
defparam memory_inst18.INIT_E = 256'h895d8501da5715979cfd60b9def311a5c23c907ba894fd50ae5bd1f3e8ed2247;
defparam memory_inst18.INIT_F = 256'h25bcdc196eb9d98bc1b5801ae65c9ce8da4b0e6d00579b309fa5041b772d47e3;

Memory memory_inst19(
    .clk(clk),
    .reset(reset),
    .addr(addr),
    .i_data_word(i_data_word),
    .o_data_byte(o_data_byte),
    .cs(cs[19]),
    .read_byte_sel(read_byte_sel),
    .rw(rw)
);
defparam memory_inst19.INIT_0 = 256'h07d9dcd9625f175da7f4ef654e89c673d8b99a55eea91cafee90f76f2d618320;
defparam memory_inst19.INIT_1 = 256'h4a740534fb1cacc2b3fa2cb3b7202aeb397a5f076d6591c6ad44476d5e347d67;
defparam memory_inst19.INIT_2 = 256'hdc1ba2d1a54e019f9d8538027a8eb47d44f29fbf5592c245d8625c78fba9ceff;
defparam memory_inst19.INIT_3 = 256'hfd9424b0769eac2c262251d471f84ce8c3b1ee61d50b5b04b06819bca53a863c;
defparam memory_inst19.INIT_4 = 256'h0a08b1e758d836b5f55bdb376c14764ff2426590752c062c1ca1dd6615d4a04d;
defparam memory_inst19.INIT_5 = 256'h117499c8db0ea1789b7db8554adc980c878be20dd6af92e8d4757ce2c6923dc7;
defparam memory_inst19.INIT_6 = 256'h7f4744ef9c5d22eba81faf26477f90f7c52e7c02613ec79c202b033b5355b4ff;
defparam memory_inst19.INIT_7 = 256'hec4e9d31fcac4ff0820f285d6b39a96afb9e4000bc1ac97b837e9431cced7f68;
defparam memory_inst19.INIT_8 = 256'h429598c3ef78e7b5e57dd1b7f7e631715ad641df8978542f84e762ec85ed8007;
defparam memory_inst19.INIT_9 = 256'h3818c9393d879df15f38a5d24c32cf78e24fe4888bf6da859adbaaf1a64f7775;
defparam memory_inst19.INIT_A = 256'h2e3267f74bca6f4cb39e16556fa95799fbcd04e80b3b45ef0f6be4208306f329;
defparam memory_inst19.INIT_B = 256'h9e228cda55f4784cf2bf72ab12569b37397cdb7c7d97309e3e0729b3050a11ef;
defparam memory_inst19.INIT_C = 256'h86ba102349ce819983688c88afcc714347d2efb058ace0bb01d51f8664d1ebd7;
defparam memory_inst19.INIT_D = 256'h720c215806df59b96471ef3cff0dc0142add109e8f3f38d43effa152a85c449a;
defparam memory_inst19.INIT_E = 256'he9fdf04f35fe0e6e15ab1636c0b1e0b1f130bef9d6e9d6ff246ed6d6c0e34841;
defparam memory_inst19.INIT_F = 256'hf9b0d206eb8041997d4b675522f6de1ef7fb15554c8e5d7fe245ea2861b608e6;


endmodule